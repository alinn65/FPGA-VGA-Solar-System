module orbit_rom_mercur (
    input wire [8:0] angle_index,  // 0-359
    output reg signed [10:0] x_out,
    output reg signed [10:0] y_out
);

always @(*) begin
    case (angle_index)
        9'd0: begin x_out = 1220; y_out = 540; end
        9'd1: begin x_out = 1219; y_out = 535; end
        9'd2: begin x_out = 1219; y_out = 530; end
        9'd3: begin x_out = 1219; y_out = 526; end
        9'd4: begin x_out = 1219; y_out = 521; end
        9'd5: begin x_out = 1219; y_out = 517; end
        9'd6: begin x_out = 1218; y_out = 512; end
        9'd7: begin x_out = 1218; y_out = 508; end
        9'd8: begin x_out = 1217; y_out = 503; end
        9'd9: begin x_out = 1216; y_out = 499; end
        9'd10: begin x_out = 1216; y_out = 494; end
        9'd11: begin x_out = 1215; y_out = 490; end
        9'd12: begin x_out = 1214; y_out = 485; end
        9'd13: begin x_out = 1213; y_out = 481; end
        9'd14: begin x_out = 1212; y_out = 477; end
        9'd15: begin x_out = 1211; y_out = 472; end
        9'd16: begin x_out = 1209; y_out = 468; end
        9'd17: begin x_out = 1208; y_out = 463; end
        9'd18: begin x_out = 1207; y_out = 459; end
        9'd19: begin x_out = 1205; y_out = 455; end
        9'd20: begin x_out = 1204; y_out = 451; end
        9'd21: begin x_out = 1202; y_out = 446; end
        9'd22: begin x_out = 1201; y_out = 442; end
        9'd23: begin x_out = 1199; y_out = 438; end
        9'd24: begin x_out = 1197; y_out = 434; end
        9'd25: begin x_out = 1195; y_out = 430; end
        9'd26: begin x_out = 1193; y_out = 426; end
        9'd27: begin x_out = 1191; y_out = 421; end
        9'd28: begin x_out = 1189; y_out = 417; end
        9'd29: begin x_out = 1187; y_out = 413; end
        9'd30: begin x_out = 1185; y_out = 410; end
        9'd31: begin x_out = 1182; y_out = 406; end
        9'd32: begin x_out = 1180; y_out = 402; end
        9'd33: begin x_out = 1178; y_out = 398; end
        9'd34: begin x_out = 1175; y_out = 394; end
        9'd35: begin x_out = 1172; y_out = 390; end
        9'd36: begin x_out = 1170; y_out = 387; end
        9'd37: begin x_out = 1167; y_out = 383; end
        9'd38: begin x_out = 1164; y_out = 379; end
        9'd39: begin x_out = 1162; y_out = 376; end
        9'd40: begin x_out = 1159; y_out = 372; end
        9'd41: begin x_out = 1156; y_out = 369; end
        9'd42: begin x_out = 1153; y_out = 366; end
        9'd43: begin x_out = 1150; y_out = 362; end
        9'd44: begin x_out = 1147; y_out = 359; end
        9'd45: begin x_out = 1143; y_out = 356; end
        9'd46: begin x_out = 1140; y_out = 352; end
        9'd47: begin x_out = 1137; y_out = 349; end
        9'd48: begin x_out = 1133; y_out = 346; end
        9'd49: begin x_out = 1130; y_out = 343; end
        9'd50: begin x_out = 1127; y_out = 340; end
        9'd51: begin x_out = 1123; y_out = 337; end
        9'd52: begin x_out = 1120; y_out = 335; end
        9'd53: begin x_out = 1116; y_out = 332; end
        9'd54: begin x_out = 1112; y_out = 329; end
        9'd55: begin x_out = 1109; y_out = 327; end
        9'd56: begin x_out = 1105; y_out = 324; end
        9'd57: begin x_out = 1101; y_out = 321; end
        9'd58: begin x_out = 1097; y_out = 319; end
        9'd59: begin x_out = 1093; y_out = 317; end
        9'd60: begin x_out = 1090; y_out = 314; end
        9'd61: begin x_out = 1086; y_out = 312; end
        9'd62: begin x_out = 1082; y_out = 310; end
        9'd63: begin x_out = 1078; y_out = 308; end
        9'd64: begin x_out = 1073; y_out = 306; end
        9'd65: begin x_out = 1069; y_out = 304; end
        9'd66: begin x_out = 1065; y_out = 302; end
        9'd67: begin x_out = 1061; y_out = 300; end
        9'd68: begin x_out = 1057; y_out = 298; end
        9'd69: begin x_out = 1053; y_out = 297; end
        9'd70: begin x_out = 1048; y_out = 295; end
        9'd71: begin x_out = 1044; y_out = 294; end
        9'd72: begin x_out = 1040; y_out = 292; end
        9'd73: begin x_out = 1036; y_out = 291; end
        9'd74: begin x_out = 1031; y_out = 290; end
        9'd75: begin x_out = 1027; y_out = 288; end
        9'd76: begin x_out = 1022; y_out = 287; end
        9'd77: begin x_out = 1018; y_out = 286; end
        9'd78: begin x_out = 1014; y_out = 285; end
        9'd79: begin x_out = 1009; y_out = 284; end
        9'd80: begin x_out = 1005; y_out = 283; end
        9'd81: begin x_out = 1000; y_out = 283; end
        9'd82: begin x_out = 996; y_out = 282; end
        9'd83: begin x_out = 991; y_out = 281; end
        9'd84: begin x_out = 987; y_out = 281; end
        9'd85: begin x_out = 982; y_out = 280; end
        9'd86: begin x_out = 978; y_out = 280; end
        9'd87: begin x_out = 973; y_out = 280; end
        9'd88: begin x_out = 969; y_out = 280; end
        9'd89: begin x_out = 964; y_out = 280; end
        9'd90: begin x_out = 960; y_out = 280; end
        9'd91: begin x_out = 955; y_out = 280; end
        9'd92: begin x_out = 950; y_out = 280; end
        9'd93: begin x_out = 946; y_out = 280; end
        9'd94: begin x_out = 941; y_out = 280; end
        9'd95: begin x_out = 937; y_out = 280; end
        9'd96: begin x_out = 932; y_out = 281; end
        9'd97: begin x_out = 928; y_out = 281; end
        9'd98: begin x_out = 923; y_out = 282; end
        9'd99: begin x_out = 919; y_out = 283; end
        9'd100: begin x_out = 914; y_out = 283; end
        9'd101: begin x_out = 910; y_out = 284; end
        9'd102: begin x_out = 905; y_out = 285; end
        9'd103: begin x_out = 901; y_out = 286; end
        9'd104: begin x_out = 897; y_out = 287; end
        9'd105: begin x_out = 892; y_out = 288; end
        9'd106: begin x_out = 888; y_out = 290; end
        9'd107: begin x_out = 883; y_out = 291; end
        9'd108: begin x_out = 879; y_out = 292; end
        9'd109: begin x_out = 875; y_out = 294; end
        9'd110: begin x_out = 871; y_out = 295; end
        9'd111: begin x_out = 866; y_out = 297; end
        9'd112: begin x_out = 862; y_out = 298; end
        9'd113: begin x_out = 858; y_out = 300; end
        9'd114: begin x_out = 854; y_out = 302; end
        9'd115: begin x_out = 850; y_out = 304; end
        9'd116: begin x_out = 846; y_out = 306; end
        9'd117: begin x_out = 841; y_out = 308; end
        9'd118: begin x_out = 837; y_out = 310; end
        9'd119: begin x_out = 833; y_out = 312; end
        9'd120: begin x_out = 830; y_out = 314; end
        9'd121: begin x_out = 826; y_out = 317; end
        9'd122: begin x_out = 822; y_out = 319; end
        9'd123: begin x_out = 818; y_out = 321; end
        9'd124: begin x_out = 814; y_out = 324; end
        9'd125: begin x_out = 810; y_out = 327; end
        9'd126: begin x_out = 807; y_out = 329; end
        9'd127: begin x_out = 803; y_out = 332; end
        9'd128: begin x_out = 799; y_out = 335; end
        9'd129: begin x_out = 796; y_out = 337; end
        9'd130: begin x_out = 792; y_out = 340; end
        9'd131: begin x_out = 789; y_out = 343; end
        9'd132: begin x_out = 786; y_out = 346; end
        9'd133: begin x_out = 782; y_out = 349; end
        9'd134: begin x_out = 779; y_out = 352; end
        9'd135: begin x_out = 776; y_out = 356; end
        9'd136: begin x_out = 772; y_out = 359; end
        9'd137: begin x_out = 769; y_out = 362; end
        9'd138: begin x_out = 766; y_out = 366; end
        9'd139: begin x_out = 763; y_out = 369; end
        9'd140: begin x_out = 760; y_out = 372; end
        9'd141: begin x_out = 757; y_out = 376; end
        9'd142: begin x_out = 755; y_out = 379; end
        9'd143: begin x_out = 752; y_out = 383; end
        9'd144: begin x_out = 749; y_out = 387; end
        9'd145: begin x_out = 747; y_out = 390; end
        9'd146: begin x_out = 744; y_out = 394; end
        9'd147: begin x_out = 741; y_out = 398; end
        9'd148: begin x_out = 739; y_out = 402; end
        9'd149: begin x_out = 737; y_out = 406; end
        9'd150: begin x_out = 734; y_out = 410; end
        9'd151: begin x_out = 732; y_out = 413; end
        9'd152: begin x_out = 730; y_out = 417; end
        9'd153: begin x_out = 728; y_out = 421; end
        9'd154: begin x_out = 726; y_out = 426; end
        9'd155: begin x_out = 724; y_out = 430; end
        9'd156: begin x_out = 722; y_out = 434; end
        9'd157: begin x_out = 720; y_out = 438; end
        9'd158: begin x_out = 718; y_out = 442; end
        9'd159: begin x_out = 717; y_out = 446; end
        9'd160: begin x_out = 715; y_out = 451; end
        9'd161: begin x_out = 714; y_out = 455; end
        9'd162: begin x_out = 712; y_out = 459; end
        9'd163: begin x_out = 711; y_out = 463; end
        9'd164: begin x_out = 710; y_out = 468; end
        9'd165: begin x_out = 708; y_out = 472; end
        9'd166: begin x_out = 707; y_out = 477; end
        9'd167: begin x_out = 706; y_out = 481; end
        9'd168: begin x_out = 705; y_out = 485; end
        9'd169: begin x_out = 704; y_out = 490; end
        9'd170: begin x_out = 703; y_out = 494; end
        9'd171: begin x_out = 703; y_out = 499; end
        9'd172: begin x_out = 702; y_out = 503; end
        9'd173: begin x_out = 701; y_out = 508; end
        9'd174: begin x_out = 701; y_out = 512; end
        9'd175: begin x_out = 700; y_out = 517; end
        9'd176: begin x_out = 700; y_out = 521; end
        9'd177: begin x_out = 700; y_out = 526; end
        9'd178: begin x_out = 700; y_out = 530; end
        9'd179: begin x_out = 700; y_out = 535; end
        9'd180: begin x_out = 700; y_out = 540; end
        9'd181: begin x_out = 700; y_out = 544; end
        9'd182: begin x_out = 700; y_out = 549; end
        9'd183: begin x_out = 700; y_out = 553; end
        9'd184: begin x_out = 700; y_out = 558; end
        9'd185: begin x_out = 700; y_out = 562; end
        9'd186: begin x_out = 701; y_out = 567; end
        9'd187: begin x_out = 701; y_out = 571; end
        9'd188: begin x_out = 702; y_out = 576; end
        9'd189: begin x_out = 703; y_out = 580; end
        9'd190: begin x_out = 703; y_out = 585; end
        9'd191: begin x_out = 704; y_out = 589; end
        9'd192: begin x_out = 705; y_out = 594; end
        9'd193: begin x_out = 706; y_out = 598; end
        9'd194: begin x_out = 707; y_out = 602; end
        9'd195: begin x_out = 708; y_out = 607; end
        9'd196: begin x_out = 710; y_out = 611; end
        9'd197: begin x_out = 711; y_out = 616; end
        9'd198: begin x_out = 712; y_out = 620; end
        9'd199: begin x_out = 714; y_out = 624; end
        9'd200: begin x_out = 715; y_out = 628; end
        9'd201: begin x_out = 717; y_out = 633; end
        9'd202: begin x_out = 718; y_out = 637; end
        9'd203: begin x_out = 720; y_out = 641; end
        9'd204: begin x_out = 722; y_out = 645; end
        9'd205: begin x_out = 724; y_out = 649; end
        9'd206: begin x_out = 726; y_out = 653; end
        9'd207: begin x_out = 728; y_out = 658; end
        9'd208: begin x_out = 730; y_out = 662; end
        9'd209: begin x_out = 732; y_out = 666; end
        9'd210: begin x_out = 734; y_out = 670; end
        9'd211: begin x_out = 737; y_out = 673; end
        9'd212: begin x_out = 739; y_out = 677; end
        9'd213: begin x_out = 741; y_out = 681; end
        9'd214: begin x_out = 744; y_out = 685; end
        9'd215: begin x_out = 747; y_out = 689; end
        9'd216: begin x_out = 749; y_out = 692; end
        9'd217: begin x_out = 752; y_out = 696; end
        9'd218: begin x_out = 755; y_out = 700; end
        9'd219: begin x_out = 757; y_out = 703; end
        9'd220: begin x_out = 760; y_out = 707; end
        9'd221: begin x_out = 763; y_out = 710; end
        9'd222: begin x_out = 766; y_out = 713; end
        9'd223: begin x_out = 769; y_out = 717; end
        9'd224: begin x_out = 772; y_out = 720; end
        9'd225: begin x_out = 776; y_out = 723; end
        9'd226: begin x_out = 779; y_out = 727; end
        9'd227: begin x_out = 782; y_out = 730; end
        9'd228: begin x_out = 786; y_out = 733; end
        9'd229: begin x_out = 789; y_out = 736; end
        9'd230: begin x_out = 792; y_out = 739; end
        9'd231: begin x_out = 796; y_out = 742; end
        9'd232: begin x_out = 799; y_out = 744; end
        9'd233: begin x_out = 803; y_out = 747; end
        9'd234: begin x_out = 807; y_out = 750; end
        9'd235: begin x_out = 810; y_out = 752; end
        9'd236: begin x_out = 814; y_out = 755; end
        9'd237: begin x_out = 818; y_out = 758; end
        9'd238: begin x_out = 822; y_out = 760; end
        9'd239: begin x_out = 826; y_out = 762; end
        9'd240: begin x_out = 829; y_out = 765; end
        9'd241: begin x_out = 833; y_out = 767; end
        9'd242: begin x_out = 837; y_out = 769; end
        9'd243: begin x_out = 841; y_out = 771; end
        9'd244: begin x_out = 846; y_out = 773; end
        9'd245: begin x_out = 850; y_out = 775; end
        9'd246: begin x_out = 854; y_out = 777; end
        9'd247: begin x_out = 858; y_out = 779; end
        9'd248: begin x_out = 862; y_out = 781; end
        9'd249: begin x_out = 866; y_out = 782; end
        9'd250: begin x_out = 871; y_out = 784; end
        9'd251: begin x_out = 875; y_out = 785; end
        9'd252: begin x_out = 879; y_out = 787; end
        9'd253: begin x_out = 883; y_out = 788; end
        9'd254: begin x_out = 888; y_out = 789; end
        9'd255: begin x_out = 892; y_out = 791; end
        9'd256: begin x_out = 897; y_out = 792; end
        9'd257: begin x_out = 901; y_out = 793; end
        9'd258: begin x_out = 905; y_out = 794; end
        9'd259: begin x_out = 910; y_out = 795; end
        9'd260: begin x_out = 914; y_out = 796; end
        9'd261: begin x_out = 919; y_out = 796; end
        9'd262: begin x_out = 923; y_out = 797; end
        9'd263: begin x_out = 928; y_out = 798; end
        9'd264: begin x_out = 932; y_out = 798; end
        9'd265: begin x_out = 937; y_out = 799; end
        9'd266: begin x_out = 941; y_out = 799; end
        9'd267: begin x_out = 946; y_out = 799; end
        9'd268: begin x_out = 950; y_out = 799; end
        9'd269: begin x_out = 955; y_out = 799; end
        9'd270: begin x_out = 960; y_out = 800; end
        9'd271: begin x_out = 964; y_out = 799; end
        9'd272: begin x_out = 969; y_out = 799; end
        9'd273: begin x_out = 973; y_out = 799; end
        9'd274: begin x_out = 978; y_out = 799; end
        9'd275: begin x_out = 982; y_out = 799; end
        9'd276: begin x_out = 987; y_out = 798; end
        9'd277: begin x_out = 991; y_out = 798; end
        9'd278: begin x_out = 996; y_out = 797; end
        9'd279: begin x_out = 1000; y_out = 796; end
        9'd280: begin x_out = 1005; y_out = 796; end
        9'd281: begin x_out = 1009; y_out = 795; end
        9'd282: begin x_out = 1014; y_out = 794; end
        9'd283: begin x_out = 1018; y_out = 793; end
        9'd284: begin x_out = 1022; y_out = 792; end
        9'd285: begin x_out = 1027; y_out = 791; end
        9'd286: begin x_out = 1031; y_out = 789; end
        9'd287: begin x_out = 1036; y_out = 788; end
        9'd288: begin x_out = 1040; y_out = 787; end
        9'd289: begin x_out = 1044; y_out = 785; end
        9'd290: begin x_out = 1048; y_out = 784; end
        9'd291: begin x_out = 1053; y_out = 782; end
        9'd292: begin x_out = 1057; y_out = 781; end
        9'd293: begin x_out = 1061; y_out = 779; end
        9'd294: begin x_out = 1065; y_out = 777; end
        9'd295: begin x_out = 1069; y_out = 775; end
        9'd296: begin x_out = 1073; y_out = 773; end
        9'd297: begin x_out = 1078; y_out = 771; end
        9'd298: begin x_out = 1082; y_out = 769; end
        9'd299: begin x_out = 1086; y_out = 767; end
        9'd300: begin x_out = 1090; y_out = 765; end
        9'd301: begin x_out = 1093; y_out = 762; end
        9'd302: begin x_out = 1097; y_out = 760; end
        9'd303: begin x_out = 1101; y_out = 758; end
        9'd304: begin x_out = 1105; y_out = 755; end
        9'd305: begin x_out = 1109; y_out = 752; end
        9'd306: begin x_out = 1112; y_out = 750; end
        9'd307: begin x_out = 1116; y_out = 747; end
        9'd308: begin x_out = 1120; y_out = 744; end
        9'd309: begin x_out = 1123; y_out = 742; end
        9'd310: begin x_out = 1127; y_out = 739; end
        9'd311: begin x_out = 1130; y_out = 736; end
        9'd312: begin x_out = 1133; y_out = 733; end
        9'd313: begin x_out = 1137; y_out = 730; end
        9'd314: begin x_out = 1140; y_out = 727; end
        9'd315: begin x_out = 1143; y_out = 723; end
        9'd316: begin x_out = 1147; y_out = 720; end
        9'd317: begin x_out = 1150; y_out = 717; end
        9'd318: begin x_out = 1153; y_out = 713; end
        9'd319: begin x_out = 1156; y_out = 710; end
        9'd320: begin x_out = 1159; y_out = 707; end
        9'd321: begin x_out = 1162; y_out = 703; end
        9'd322: begin x_out = 1164; y_out = 700; end
        9'd323: begin x_out = 1167; y_out = 696; end
        9'd324: begin x_out = 1170; y_out = 692; end
        9'd325: begin x_out = 1172; y_out = 689; end
        9'd326: begin x_out = 1175; y_out = 685; end
        9'd327: begin x_out = 1178; y_out = 681; end
        9'd328: begin x_out = 1180; y_out = 677; end
        9'd329: begin x_out = 1182; y_out = 673; end
        9'd330: begin x_out = 1185; y_out = 670; end
        9'd331: begin x_out = 1187; y_out = 666; end
        9'd332: begin x_out = 1189; y_out = 662; end
        9'd333: begin x_out = 1191; y_out = 658; end
        9'd334: begin x_out = 1193; y_out = 653; end
        9'd335: begin x_out = 1195; y_out = 649; end
        9'd336: begin x_out = 1197; y_out = 645; end
        9'd337: begin x_out = 1199; y_out = 641; end
        9'd338: begin x_out = 1201; y_out = 637; end
        9'd339: begin x_out = 1202; y_out = 633; end
        9'd340: begin x_out = 1204; y_out = 628; end
        9'd341: begin x_out = 1205; y_out = 624; end
        9'd342: begin x_out = 1207; y_out = 620; end
        9'd343: begin x_out = 1208; y_out = 616; end
        9'd344: begin x_out = 1209; y_out = 611; end
        9'd345: begin x_out = 1211; y_out = 607; end
        9'd346: begin x_out = 1212; y_out = 602; end
        9'd347: begin x_out = 1213; y_out = 598; end
        9'd348: begin x_out = 1214; y_out = 594; end
        9'd349: begin x_out = 1215; y_out = 589; end
        9'd350: begin x_out = 1216; y_out = 585; end
        9'd351: begin x_out = 1216; y_out = 580; end
        9'd352: begin x_out = 1217; y_out = 576; end
        9'd353: begin x_out = 1218; y_out = 571; end
        9'd354: begin x_out = 1218; y_out = 567; end
        9'd355: begin x_out = 1219; y_out = 562; end
        9'd356: begin x_out = 1219; y_out = 558; end
        9'd357: begin x_out = 1219; y_out = 553; end
        9'd358: begin x_out = 1219; y_out = 549; end

        default: begin x_out = 0; y_out = 0; end
    endcase
end

endmodule