module orbit_rom_venus (
    input wire [8:0] angle_index,  // 0-359
    output reg signed [10:0] x_out,
    output reg signed [10:0] y_out
);

always @(*) begin
    case (angle_index)
        9'd0: begin x_out = 1340; y_out = 540; end
        9'd1: begin x_out = 1339; y_out = 533; end
        9'd2: begin x_out = 1339; y_out = 526; end
        9'd3: begin x_out = 1339; y_out = 520; end
        9'd4: begin x_out = 1339; y_out = 513; end
        9'd5: begin x_out = 1338; y_out = 506; end
        9'd6: begin x_out = 1337; y_out = 500; end
        9'd7: begin x_out = 1337; y_out = 493; end
        9'd8: begin x_out = 1336; y_out = 487; end
        9'd9: begin x_out = 1335; y_out = 480; end
        9'd10: begin x_out = 1334; y_out = 474; end
        9'd11: begin x_out = 1333; y_out = 467; end
        9'd12: begin x_out = 1331; y_out = 460; end
        9'd13: begin x_out = 1330; y_out = 454; end
        9'd14: begin x_out = 1328; y_out = 448; end
        9'd15: begin x_out = 1327; y_out = 441; end
        9'd16: begin x_out = 1325; y_out = 435; end
        9'd17: begin x_out = 1323; y_out = 428; end
        9'd18: begin x_out = 1321; y_out = 422; end
        9'd19: begin x_out = 1319; y_out = 416; end
        9'd20: begin x_out = 1317; y_out = 410; end
        9'd21: begin x_out = 1314; y_out = 403; end
        9'd22: begin x_out = 1312; y_out = 397; end
        9'd23: begin x_out = 1309; y_out = 391; end
        9'd24: begin x_out = 1307; y_out = 385; end
        9'd25: begin x_out = 1304; y_out = 379; end
        9'd26: begin x_out = 1301; y_out = 373; end
        9'd27: begin x_out = 1298; y_out = 367; end
        9'd28: begin x_out = 1295; y_out = 361; end
        9'd29: begin x_out = 1292; y_out = 355; end
        9'd30: begin x_out = 1289; y_out = 350; end
        9'd31: begin x_out = 1285; y_out = 344; end
        9'd32: begin x_out = 1282; y_out = 338; end
        9'd33: begin x_out = 1278; y_out = 333; end
        9'd34: begin x_out = 1275; y_out = 327; end
        9'd35: begin x_out = 1271; y_out = 322; end
        9'd36: begin x_out = 1267; y_out = 316; end
        9'd37: begin x_out = 1263; y_out = 311; end
        9'd38: begin x_out = 1259; y_out = 306; end
        9'd39: begin x_out = 1255; y_out = 300; end
        9'd40: begin x_out = 1251; y_out = 295; end
        9'd41: begin x_out = 1246; y_out = 290; end
        9'd42: begin x_out = 1242; y_out = 285; end
        9'd43: begin x_out = 1237; y_out = 280; end
        9'd44: begin x_out = 1233; y_out = 276; end
        9'd45: begin x_out = 1228; y_out = 271; end
        9'd46: begin x_out = 1223; y_out = 266; end
        9'd47: begin x_out = 1219; y_out = 262; end
        9'd48: begin x_out = 1214; y_out = 257; end
        9'd49: begin x_out = 1209; y_out = 253; end
        9'd50: begin x_out = 1204; y_out = 248; end
        9'd51: begin x_out = 1199; y_out = 244; end
        9'd52: begin x_out = 1193; y_out = 240; end
        9'd53: begin x_out = 1188; y_out = 236; end
        9'd54: begin x_out = 1183; y_out = 232; end
        9'd55: begin x_out = 1177; y_out = 228; end
        9'd56: begin x_out = 1172; y_out = 224; end
        9'd57: begin x_out = 1166; y_out = 221; end
        9'd58: begin x_out = 1161; y_out = 217; end
        9'd59: begin x_out = 1155; y_out = 214; end
        9'd60: begin x_out = 1150; y_out = 210; end
        9'd61: begin x_out = 1144; y_out = 207; end
        9'd62: begin x_out = 1138; y_out = 204; end
        9'd63: begin x_out = 1132; y_out = 201; end
        9'd64: begin x_out = 1126; y_out = 198; end
        9'd65: begin x_out = 1120; y_out = 195; end
        9'd66: begin x_out = 1114; y_out = 192; end
        9'd67: begin x_out = 1108; y_out = 190; end
        9'd68: begin x_out = 1102; y_out = 187; end
        9'd69: begin x_out = 1096; y_out = 185; end
        9'd70: begin x_out = 1089; y_out = 182; end
        9'd71: begin x_out = 1083; y_out = 180; end
        9'd72: begin x_out = 1077; y_out = 178; end
        9'd73: begin x_out = 1071; y_out = 176; end
        9'd74: begin x_out = 1064; y_out = 174; end
        9'd75: begin x_out = 1058; y_out = 172; end
        9'd76: begin x_out = 1051; y_out = 171; end
        9'd77: begin x_out = 1045; y_out = 169; end
        9'd78: begin x_out = 1039; y_out = 168; end
        9'd79: begin x_out = 1032; y_out = 166; end
        9'd80: begin x_out = 1025; y_out = 165; end
        9'd81: begin x_out = 1019; y_out = 164; end
        9'd82: begin x_out = 1012; y_out = 163; end
        9'd83: begin x_out = 1006; y_out = 162; end
        9'd84: begin x_out = 999; y_out = 162; end
        9'd85: begin x_out = 993; y_out = 161; end
        9'd86: begin x_out = 986; y_out = 160; end
        9'd87: begin x_out = 979; y_out = 160; end
        9'd88: begin x_out = 973; y_out = 160; end
        9'd89: begin x_out = 966; y_out = 160; end
        9'd90: begin x_out = 960; y_out = 160; end
        9'd91: begin x_out = 953; y_out = 160; end
        9'd92: begin x_out = 946; y_out = 160; end
        9'd93: begin x_out = 940; y_out = 160; end
        9'd94: begin x_out = 933; y_out = 160; end
        9'd95: begin x_out = 926; y_out = 161; end
        9'd96: begin x_out = 920; y_out = 162; end
        9'd97: begin x_out = 913; y_out = 162; end
        9'd98: begin x_out = 907; y_out = 163; end
        9'd99: begin x_out = 900; y_out = 164; end
        9'd100: begin x_out = 894; y_out = 165; end
        9'd101: begin x_out = 887; y_out = 166; end
        9'd102: begin x_out = 880; y_out = 168; end
        9'd103: begin x_out = 874; y_out = 169; end
        9'd104: begin x_out = 868; y_out = 171; end
        9'd105: begin x_out = 861; y_out = 172; end
        9'd106: begin x_out = 855; y_out = 174; end
        9'd107: begin x_out = 848; y_out = 176; end
        9'd108: begin x_out = 842; y_out = 178; end
        9'd109: begin x_out = 836; y_out = 180; end
        9'd110: begin x_out = 830; y_out = 182; end
        9'd111: begin x_out = 823; y_out = 185; end
        9'd112: begin x_out = 817; y_out = 187; end
        9'd113: begin x_out = 811; y_out = 190; end
        9'd114: begin x_out = 805; y_out = 192; end
        9'd115: begin x_out = 799; y_out = 195; end
        9'd116: begin x_out = 793; y_out = 198; end
        9'd117: begin x_out = 787; y_out = 201; end
        9'd118: begin x_out = 781; y_out = 204; end
        9'd119: begin x_out = 775; y_out = 207; end
        9'd120: begin x_out = 770; y_out = 210; end
        9'd121: begin x_out = 764; y_out = 214; end
        9'd122: begin x_out = 758; y_out = 217; end
        9'd123: begin x_out = 753; y_out = 221; end
        9'd124: begin x_out = 747; y_out = 224; end
        9'd125: begin x_out = 742; y_out = 228; end
        9'd126: begin x_out = 736; y_out = 232; end
        9'd127: begin x_out = 731; y_out = 236; end
        9'd128: begin x_out = 726; y_out = 240; end
        9'd129: begin x_out = 720; y_out = 244; end
        9'd130: begin x_out = 715; y_out = 248; end
        9'd131: begin x_out = 710; y_out = 253; end
        9'd132: begin x_out = 705; y_out = 257; end
        9'd133: begin x_out = 700; y_out = 262; end
        9'd134: begin x_out = 696; y_out = 266; end
        9'd135: begin x_out = 691; y_out = 271; end
        9'd136: begin x_out = 686; y_out = 276; end
        9'd137: begin x_out = 682; y_out = 280; end
        9'd138: begin x_out = 677; y_out = 285; end
        9'd139: begin x_out = 673; y_out = 290; end
        9'd140: begin x_out = 668; y_out = 295; end
        9'd141: begin x_out = 664; y_out = 300; end
        9'd142: begin x_out = 660; y_out = 306; end
        9'd143: begin x_out = 656; y_out = 311; end
        9'd144: begin x_out = 652; y_out = 316; end
        9'd145: begin x_out = 648; y_out = 322; end
        9'd146: begin x_out = 644; y_out = 327; end
        9'd147: begin x_out = 641; y_out = 333; end
        9'd148: begin x_out = 637; y_out = 338; end
        9'd149: begin x_out = 634; y_out = 344; end
        9'd150: begin x_out = 630; y_out = 350; end
        9'd151: begin x_out = 627; y_out = 355; end
        9'd152: begin x_out = 624; y_out = 361; end
        9'd153: begin x_out = 621; y_out = 367; end
        9'd154: begin x_out = 618; y_out = 373; end
        9'd155: begin x_out = 615; y_out = 379; end
        9'd156: begin x_out = 612; y_out = 385; end
        9'd157: begin x_out = 610; y_out = 391; end
        9'd158: begin x_out = 607; y_out = 397; end
        9'd159: begin x_out = 605; y_out = 403; end
        9'd160: begin x_out = 602; y_out = 410; end
        9'd161: begin x_out = 600; y_out = 416; end
        9'd162: begin x_out = 598; y_out = 422; end
        9'd163: begin x_out = 596; y_out = 428; end
        9'd164: begin x_out = 594; y_out = 435; end
        9'd165: begin x_out = 592; y_out = 441; end
        9'd166: begin x_out = 591; y_out = 448; end
        9'd167: begin x_out = 589; y_out = 454; end
        9'd168: begin x_out = 588; y_out = 460; end
        9'd169: begin x_out = 586; y_out = 467; end
        9'd170: begin x_out = 585; y_out = 474; end
        9'd171: begin x_out = 584; y_out = 480; end
        9'd172: begin x_out = 583; y_out = 487; end
        9'd173: begin x_out = 582; y_out = 493; end
        9'd174: begin x_out = 582; y_out = 500; end
        9'd175: begin x_out = 581; y_out = 506; end
        9'd176: begin x_out = 580; y_out = 513; end
        9'd177: begin x_out = 580; y_out = 520; end
        9'd178: begin x_out = 580; y_out = 526; end
        9'd179: begin x_out = 580; y_out = 533; end
        9'd180: begin x_out = 580; y_out = 540; end
        9'd181: begin x_out = 580; y_out = 546; end
        9'd182: begin x_out = 580; y_out = 553; end
        9'd183: begin x_out = 580; y_out = 559; end
        9'd184: begin x_out = 580; y_out = 566; end
        9'd185: begin x_out = 581; y_out = 573; end
        9'd186: begin x_out = 582; y_out = 579; end
        9'd187: begin x_out = 582; y_out = 586; end
        9'd188: begin x_out = 583; y_out = 592; end
        9'd189: begin x_out = 584; y_out = 599; end
        9'd190: begin x_out = 585; y_out = 605; end
        9'd191: begin x_out = 586; y_out = 612; end
        9'd192: begin x_out = 588; y_out = 619; end
        9'd193: begin x_out = 589; y_out = 625; end
        9'd194: begin x_out = 591; y_out = 631; end
        9'd195: begin x_out = 592; y_out = 638; end
        9'd196: begin x_out = 594; y_out = 644; end
        9'd197: begin x_out = 596; y_out = 651; end
        9'd198: begin x_out = 598; y_out = 657; end
        9'd199: begin x_out = 600; y_out = 663; end
        9'd200: begin x_out = 602; y_out = 669; end
        9'd201: begin x_out = 605; y_out = 676; end
        9'd202: begin x_out = 607; y_out = 682; end
        9'd203: begin x_out = 610; y_out = 688; end
        9'd204: begin x_out = 612; y_out = 694; end
        9'd205: begin x_out = 615; y_out = 700; end
        9'd206: begin x_out = 618; y_out = 706; end
        9'd207: begin x_out = 621; y_out = 712; end
        9'd208: begin x_out = 624; y_out = 718; end
        9'd209: begin x_out = 627; y_out = 724; end
        9'd210: begin x_out = 630; y_out = 730; end
        9'd211: begin x_out = 634; y_out = 735; end
        9'd212: begin x_out = 637; y_out = 741; end
        9'd213: begin x_out = 641; y_out = 746; end
        9'd214: begin x_out = 644; y_out = 752; end
        9'd215: begin x_out = 648; y_out = 757; end
        9'd216: begin x_out = 652; y_out = 763; end
        9'd217: begin x_out = 656; y_out = 768; end
        9'd218: begin x_out = 660; y_out = 773; end
        9'd219: begin x_out = 664; y_out = 779; end
        9'd220: begin x_out = 668; y_out = 784; end
        9'd221: begin x_out = 673; y_out = 789; end
        9'd222: begin x_out = 677; y_out = 794; end
        9'd223: begin x_out = 682; y_out = 799; end
        9'd224: begin x_out = 686; y_out = 803; end
        9'd225: begin x_out = 691; y_out = 808; end
        9'd226: begin x_out = 696; y_out = 813; end
        9'd227: begin x_out = 700; y_out = 817; end
        9'd228: begin x_out = 705; y_out = 822; end
        9'd229: begin x_out = 710; y_out = 826; end
        9'd230: begin x_out = 715; y_out = 831; end
        9'd231: begin x_out = 720; y_out = 835; end
        9'd232: begin x_out = 726; y_out = 839; end
        9'd233: begin x_out = 731; y_out = 843; end
        9'd234: begin x_out = 736; y_out = 847; end
        9'd235: begin x_out = 742; y_out = 851; end
        9'd236: begin x_out = 747; y_out = 855; end
        9'd237: begin x_out = 753; y_out = 858; end
        9'd238: begin x_out = 758; y_out = 862; end
        9'd239: begin x_out = 764; y_out = 865; end
        9'd240: begin x_out = 769; y_out = 869; end
        9'd241: begin x_out = 775; y_out = 872; end
        9'd242: begin x_out = 781; y_out = 875; end
        9'd243: begin x_out = 787; y_out = 878; end
        9'd244: begin x_out = 793; y_out = 881; end
        9'd245: begin x_out = 799; y_out = 884; end
        9'd246: begin x_out = 805; y_out = 887; end
        9'd247: begin x_out = 811; y_out = 889; end
        9'd248: begin x_out = 817; y_out = 892; end
        9'd249: begin x_out = 823; y_out = 894; end
        9'd250: begin x_out = 830; y_out = 897; end
        9'd251: begin x_out = 836; y_out = 899; end
        9'd252: begin x_out = 842; y_out = 901; end
        9'd253: begin x_out = 848; y_out = 903; end
        9'd254: begin x_out = 855; y_out = 905; end
        9'd255: begin x_out = 861; y_out = 907; end
        9'd256: begin x_out = 868; y_out = 908; end
        9'd257: begin x_out = 874; y_out = 910; end
        9'd258: begin x_out = 880; y_out = 911; end
        9'd259: begin x_out = 887; y_out = 913; end
        9'd260: begin x_out = 894; y_out = 914; end
        9'd261: begin x_out = 900; y_out = 915; end
        9'd262: begin x_out = 907; y_out = 916; end
        9'd263: begin x_out = 913; y_out = 917; end
        9'd264: begin x_out = 920; y_out = 917; end
        9'd265: begin x_out = 926; y_out = 918; end
        9'd266: begin x_out = 933; y_out = 919; end
        9'd267: begin x_out = 940; y_out = 919; end
        9'd268: begin x_out = 946; y_out = 919; end
        9'd269: begin x_out = 953; y_out = 919; end
        9'd270: begin x_out = 959; y_out = 920; end
        9'd271: begin x_out = 966; y_out = 919; end
        9'd272: begin x_out = 973; y_out = 919; end
        9'd273: begin x_out = 979; y_out = 919; end
        9'd274: begin x_out = 986; y_out = 919; end
        9'd275: begin x_out = 993; y_out = 918; end
        9'd276: begin x_out = 999; y_out = 917; end
        9'd277: begin x_out = 1006; y_out = 917; end
        9'd278: begin x_out = 1012; y_out = 916; end
        9'd279: begin x_out = 1019; y_out = 915; end
        9'd280: begin x_out = 1025; y_out = 914; end
        9'd281: begin x_out = 1032; y_out = 913; end
        9'd282: begin x_out = 1039; y_out = 911; end
        9'd283: begin x_out = 1045; y_out = 910; end
        9'd284: begin x_out = 1051; y_out = 908; end
        9'd285: begin x_out = 1058; y_out = 907; end
        9'd286: begin x_out = 1064; y_out = 905; end
        9'd287: begin x_out = 1071; y_out = 903; end
        9'd288: begin x_out = 1077; y_out = 901; end
        9'd289: begin x_out = 1083; y_out = 899; end
        9'd290: begin x_out = 1089; y_out = 897; end
        9'd291: begin x_out = 1096; y_out = 894; end
        9'd292: begin x_out = 1102; y_out = 892; end
        9'd293: begin x_out = 1108; y_out = 889; end
        9'd294: begin x_out = 1114; y_out = 887; end
        9'd295: begin x_out = 1120; y_out = 884; end
        9'd296: begin x_out = 1126; y_out = 881; end
        9'd297: begin x_out = 1132; y_out = 878; end
        9'd298: begin x_out = 1138; y_out = 875; end
        9'd299: begin x_out = 1144; y_out = 872; end
        9'd300: begin x_out = 1150; y_out = 869; end
        9'd301: begin x_out = 1155; y_out = 865; end
        9'd302: begin x_out = 1161; y_out = 862; end
        9'd303: begin x_out = 1166; y_out = 858; end
        9'd304: begin x_out = 1172; y_out = 855; end
        9'd305: begin x_out = 1177; y_out = 851; end
        9'd306: begin x_out = 1183; y_out = 847; end
        9'd307: begin x_out = 1188; y_out = 843; end
        9'd308: begin x_out = 1193; y_out = 839; end
        9'd309: begin x_out = 1199; y_out = 835; end
        9'd310: begin x_out = 1204; y_out = 831; end
        9'd311: begin x_out = 1209; y_out = 826; end
        9'd312: begin x_out = 1214; y_out = 822; end
        9'd313: begin x_out = 1219; y_out = 817; end
        9'd314: begin x_out = 1223; y_out = 813; end
        9'd315: begin x_out = 1228; y_out = 808; end
        9'd316: begin x_out = 1233; y_out = 803; end
        9'd317: begin x_out = 1237; y_out = 799; end
        9'd318: begin x_out = 1242; y_out = 794; end
        9'd319: begin x_out = 1246; y_out = 789; end
        9'd320: begin x_out = 1251; y_out = 784; end
        9'd321: begin x_out = 1255; y_out = 779; end
        9'd322: begin x_out = 1259; y_out = 773; end
        9'd323: begin x_out = 1263; y_out = 768; end
        9'd324: begin x_out = 1267; y_out = 763; end
        9'd325: begin x_out = 1271; y_out = 757; end
        9'd326: begin x_out = 1275; y_out = 752; end
        9'd327: begin x_out = 1278; y_out = 746; end
        9'd328: begin x_out = 1282; y_out = 741; end
        9'd329: begin x_out = 1285; y_out = 735; end
        9'd330: begin x_out = 1289; y_out = 730; end
        9'd331: begin x_out = 1292; y_out = 724; end
        9'd332: begin x_out = 1295; y_out = 718; end
        9'd333: begin x_out = 1298; y_out = 712; end
        9'd334: begin x_out = 1301; y_out = 706; end
        9'd335: begin x_out = 1304; y_out = 700; end
        9'd336: begin x_out = 1307; y_out = 694; end
        9'd337: begin x_out = 1309; y_out = 688; end
        9'd338: begin x_out = 1312; y_out = 682; end
        9'd339: begin x_out = 1314; y_out = 676; end
        9'd340: begin x_out = 1317; y_out = 669; end
        9'd341: begin x_out = 1319; y_out = 663; end
        9'd342: begin x_out = 1321; y_out = 657; end
        9'd343: begin x_out = 1323; y_out = 651; end
        9'd344: begin x_out = 1325; y_out = 644; end
        9'd345: begin x_out = 1327; y_out = 638; end
        9'd346: begin x_out = 1328; y_out = 631; end
        9'd347: begin x_out = 1330; y_out = 625; end
        9'd348: begin x_out = 1331; y_out = 619; end
        9'd349: begin x_out = 1333; y_out = 612; end
        9'd350: begin x_out = 1334; y_out = 605; end
        9'd351: begin x_out = 1335; y_out = 599; end
        9'd352: begin x_out = 1336; y_out = 592; end
        9'd353: begin x_out = 1337; y_out = 586; end
        9'd354: begin x_out = 1337; y_out = 579; end
        9'd355: begin x_out = 1338; y_out = 573; end
        9'd356: begin x_out = 1339; y_out = 566; end
        9'd357: begin x_out = 1339; y_out = 559; end
        9'd358: begin x_out = 1339; y_out = 553; end

        default: begin x_out = 0; y_out = 0; end
    endcase
end

endmodule